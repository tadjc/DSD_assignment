module BUFFER(out, in);
input in;
output out;

assign out = in;
endmodule