module dtat_path_test_1()
endmodule